.subckt IDEAL_INVERTER in out vdd vss
B_INV out vss V = V(in) > V(vdd)/2 ? V(vss) : V(vdd)
.ENDS