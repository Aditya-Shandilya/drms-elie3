.subckt Ideal_inv in out vdd vss
B_INV out vss V = V(in) > V(vdd)/2 ? V(vss) : V(vdd)
.ends Ideal_inv