* Ideal Decimator

.subckt ideal_decimator analog_in analog_clk adaclout adaccout samples=512

*Input Interface
abridge_in [analog_in] [din] adc_buff
abridge_clk [analog_clk] [dclk] adc_buff
.model adc_buff adc_bridge(in_low = 1.5 in_high = 1.5)
ainv din dinb inv_gate
.model inv_gate d_inverter(rise_delay = 1e-9 fall_delay = 1e-9)

*The Counter (Accumulator)
XCounter din dinb dclk dreset dout1 dout2 dout3 dout4 dout5 dout6 dout7 dout8 dout9 dout10 count10

*The Latch (Sample & Hold)
Xlatch dout1 dout2 dout3 dout4 dout5 dout6 dout7 dout8 dout9 dout10
+ dlout1 dlout2 dlout3 dlout4 dlout5 dlout6 dlout7 dlout8 dlout9 dlout10 dlatch_clk
+ latch10

*Control Logic
adivn dclk ddivn divider
.model divider d_fdiv(div_factor = 'samples' high_cycles = 1
+ i_count = 0 rise_delay = 1e-9 fall_delay = 1e-9)
adelay1 ddivn dlatch_clk buff_delay
adelay2 dlatch_clk dreset buff_delay
.model buff_delay d_buffer(rise_delay = 10n fall_delay = 10n input_load = 0.5e-12)

*DAC 1: Latched Output (The Stepped Sine Wave)
Xdac_latch dlout1 dlout2 dlout3 dlout4 dlout5 dlout6 dlout7 dlout8 dlout9 dlout10 adaclout dac10

*DAC 2: Real-time Counter (The Blue Sawtooth)
Xdac_counter dout1 dout2 dout3 dout4 dout5 dout6 dout7 dout8 dout9 dout10 adaccout dac10

*Load dependencies
.include count-latch-dac.cir

.ends ideal_decimator